`timescale 1ns / 1ps

module memory(
    input wire clk,        // сигнал синхронизации
    input wire WE,         // сигнал разрешения записи данных
    input wire [31:0] A,   // адрес данных для чтения или записи данных
    input wire [31:0] WD,  // данные для записи
    output reg [31:0] RD = 0   // прочитанные данные
);
    
reg [31:0] RAM [0:127]; // 128 регистров, каждый из которых имеет разрядность в 32 бита
integer i = 0;
 
// инициализируем память нулями
initial
begin
   for(i = 0;i<128;i++)
   begin
       RAM[i] = 0;
   end
end

always @(posedge clk)
begin
   if(WE) // если активен сигнал разрешения записи данных, то начинаем записывать данные
    begin
        RAM[A[31:2]] <= WD; // вместо того, чтобы считвать 1 байт, считываем целое слово
    end
   
   else // если неактивен сигнал разрешения записи, то производится считывание данных из памяти
    begin
       RD <= RAM[A[31:2]];  
    end 
end

endmodule
